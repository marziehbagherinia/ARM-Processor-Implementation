library verilog;
use verilog.vl_types.all;
entity InstructionMemory is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        address         : in     vl_logic_vector(31 downto 0);
        WriteData       : in     vl_logic_vector(31 downto 0);
        MemRead         : in     vl_logic;
        MemWrite        : in     vl_logic;
        ReadData        : out    vl_logic_vector(31 downto 0)
    );
end InstructionMemory;
